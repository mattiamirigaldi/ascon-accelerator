package ascon_pkg;
  typedef logic [4:0][63:0] state_t;
endpackage : ascon_pkg
